----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:51:15 10/18/2022 
-- Design Name: 
-- Module Name:    Control_Unit - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;




-- if load word or store word then ALU op <= Add instruction .

entity Control_Unit is
	Port ( 
				Op_code : in std_logic_vector ( 5 downto 0 ) ;

				PC_src : out std_logic;

				ALU_Src : out std_logic;
				Mem_write :out std_logic;
				Reg_write :out std_logic;
				Reg_dst :out std_logic;
				ALU_op : out std_logic_vector( 1 downto 0 ) ;
				Mem_to_reg : out std_logic;
				Mem_read : out std_logic;
				Branch : out std_logic
				);
end Control_Unit;

architecture Behavioral of Control_Unit is

begin
	process(clk,op_code)
		begin 
			if(clk_rising) then 
				case Op_code is
					when "000000" =>
					-- depends on function code 
						ALU_op<="10";
						Reg_dst<='1';
						ALU_Src<='0';
						Reg_write<'1';
						Mem_write<='0';
						Mem_read<='0';
						Mem_to_reg<='0';
					when "100011" =>
					-- load word
					
					when "101011" =>
					-- store word 
					
					-------------------------------------
					----- I type instructions ------------------
					when "001001" =>
					-- add imm
					
					when "001010" =>
					--set less than imm
					
					when "001011" =>
					--set less than imm unsigned
					
					when "001100" =>
					-- AND imm
					
					when "001101" =>
					-- OR imm 
					
					when "001110" =>
					--XOR immediate
					
					-------------------------------------------
					----- jump instrucions --------------------
					
				
				end case;
		
		
		
			end if;
		end process;


end Behavioral;

